FULL_CIR_SIM
**********************************************************************************************************
* SOLAR MAX. POWER POINT TRACKER MQP
* JOHNATHAN ADAMS, BENJAMIN BEAUREGARD, ANDREW FLYNN
* ADVISOR: PROFESSOR ALEXANDER EMANUEL
* A, B, C TERM 2016-2017
* WORCESTER POLYTECHNIC INSTITUTE
**********************************************************************************************************
* DOCUMENT: FULL_CIR_SIM.CIR
* DATE CREATED: 10/12/16

**********************************************************************************************************
* INCLUDE: LIBRARY AND EXTERNAL FILE INCLUDES
**********************************************************************************************************
.LIB MPPT_MODELS.LIB

**********************************************************************************************************
* MAIN: FOR CONNECTING PRIMARY SUBCIRCUITS TOGETHER
**********************************************************************************************************
XSOLAR 1 0 SOLAR_SIM
*VTEST 1 0 30
XFILTER_1 1 2 0 FILTER_1
*.OPTIONS <Parameter Name>={SCHEDULE(<time-value>, <parameter value>
.PARAM WIDTH=0.01m
VPWM1 3 4 PULSE(0 3.3 0 500n 500n {WIDTH} 0.02m)
XMPPT_BUCK 2 3 4 5 0 MPPT_BUCK
*XFILTER_2 5 6 0 FILTER_2
*VPWM2 7 8 PULSE(0 3.3 0 1n 1n 0.01m 0.02m)
*XOUT_BUCK 6 7 8 9 0 OUT_BUCK
RLOAD 5 0 100

**********************************************************************************************************
* SOLAR CELL SIMULATOR
* OUTPUT NODES TO BE CONNECTED TO FILTER
* GND_REF TO BE CONNECTED TO NODE 0
**********************************************************************************************************
.SUBCKT SOLAR_SIM P_OUT GND
    VSOLAR 2 1 30
    D1 2 P_OUT D1N4004
    RSOLAR1 P_OUT 3 10K
    * RSOLAR1 AND RSOLAR2 MAKE UP 50% 10K POT TO IRF1310 GATE
    RSOLAR2 3 4 5K
    RSOLAR3 4 1 5K
    XQ1 GND 4 1 IRF1310
.ENDS
* END SOLAR_SIM

**********************************************************************************************************
* FILTER 1
* INPUT NODES TO BE CONNECTED TO SOLAR CELL SIMULATOR OUTPUT
* OUTPUT NODES TO BE CONNECTED TO BUCK CONVERTER INPUT
**********************************************************************************************************
.SUBCKT FILTER_1 P_IN P_OUT GND
	XFLTR1 P_IN 1 GND FLTR_STAGE
	XFLTR2 1 2 GND FLTR_STAGE
	LFLTR_FINAL 2 3 1m
	RIND_FLTR_FINAL 3 P_OUT 10m
	CFLTR_FINAL 4 GND 33n
	RCAP_FLTR_FINAL P_OUT 4 8m
	D_FREE P_OUT P_IN MBR1060
	LOUT_FLTR P_REF 1 1m
	RIND_OUT_FLTR 1 P_OUT 137m
	COUT_FLTR 2 GND 15u
	RCAP_OUT_FLTR P_OUT 2 8m
.ENDS
*END FILTER_1

.SUBCKT FLTR_STAGE 1 2 3
    * External node designations:
    * Node 1 -> stage input
    * Node 2 -> stage output
    * Node 3 -> ground
    L 1 4 1m
    R_IND 4 2 10m
    C 5 3 100n
    R_CAP 5 2 8m
.ENDS
* END FLTR_STAGE

**********************************************************************************************************
* MPPT BUCK CONVERTER
* INPUT NODES TO BE CONNECTED TO FILTER OUTPUT
* SIG_IN NODE TO BE CONNECTED TO PULSE VOLTAGE SOURCE IN MAIN FOR PWM
* OUTPUT NODES TO BE CONNECTED TO FILTER 2
**********************************************************************************************************
.SUBCKT MPPT_BUCK P_IN SIG_IN P_REF P_OUT GND
	XQ2 P_IN SIG_IN P_REF DMT6009LCT
	D2 GND P_REF MBR1060
	LOUT_FLTR P_REF 1 1m
	RIND_OUT_FLTR 1 P_OUT 137m
	COUT_FLTR 2 GND 15u
	RCAP_OUT_FLTR P_OUT 2 8m
.ENDS
* END MPPT_BUCK

**********************************************************************************************************
* FILTER 2
* INPUT NODES TO BE CONNECTED TO MPPT BUCK CONVERTER OUTPUT
* OUTPUT NODES TO BE CONNECTED TO OUTPUT BUCK CONVERTER INPUT
* NOTE: USES "FLTR_STAGE" SUBCIRCUIT FROM FILTER 1
**********************************************************************************************************
.SUBCKT FILTER_2 P_IN P_OUT GND
	XFLTR1 P_IN 1 GND FLTR_STAGE
	XFLTR2 1 2 GND FLTR_STAGE
	LFLTR_FINAL 2 3 1m
	RIND_FLTR_FINAL 3 P_OUT 10m
	CFLTR_FINAL 4 GND 33n
	RCAP_FLTR_FINAL P_OUT 4 8m
	D_FREE P_OUT P_IN MBR1060
	LOUT_FLTR P_REF 1 1m
	RIND_OUT_FLTR 1 P_OUT 137m
	COUT_FLTR 2 GND 15u
	RCAP_OUT_FLTR P_OUT 2 8m
.ENDS
*END FILTER_2

**********************************************************************************************************
* OUT BUCK CONVERTER
* P_IN AND GND NODES TO BE CONNECTED TO FILTER_2 OUTPUT
* SIG_IN NODE TO BE CONNECTED TO PULSE VOLTAGE SOURCE IN MAIN FOR PWM
* OUTPUT NODES TO BE CONNECTED TO LOAD (IN MAIN)
* NOTE: USES DMT6009LCT SUBCIRCUIT FROM MPPT_BUCK
**********************************************************************************************************
.SUBCKT OUT_BUCK P_IN SIG_IN P_REF P_OUT GND
	XQ3 P_IN SIG_IN P_REF DMT6009LCT
	D3 GND P_REF MBR1060
	LOUT_FLTR P_REF 1 1m
	RIND_OUT_FLTR 1 P_OUT 137m
	COUT_FLTR 2 GND 15u
	RCAP_OUT_FLTR P_OUT 2 8m
.ENDS
* END OUT_BUCK

**********************************************************************************************************
* SIMULATION CONFIGURATION
**********************************************************************************************************
.PROBE
.TRAN 50m 50m 0u 1u UIC
*.DC PARAM WIDTH LIST 0.005m 0.01m 0.015m
.END 

PWM_TRIAL_320
.LIB BRUTE_FORCE_VOLTAGE_SOURCE.LIB
XV1 1 0 PWM
.PROBE
.TRAN 1580m 1580m 0u 1u UIC
.END
PWM_TRIAL_2
*
* INPUT VOLTAGE
VIN	1	0	SIN(5V 4V 500HZ)    ;SIN(VOffset VPeak Frequency)
RIN	1	0	1K
*
* 10KHZ TRIANGLE WAVE 
* (GENERATED USING PULSE SOURCE WITH LONG RISE/FALL TIMES)
VTRI	2	0	PULSE(0V 10V 0 49US 49US 1US 100US)
RTRI	2	0	1MEG
*
* COMPARATOR, INPUT = V(1,2)
* FOR V(1,2) < -1MV, OUTPUT = 0V
* FOR V(1,2) > +1MV, OUTPUT = 10V
ECOMP	3	0	TABLE {V(1,2)} = (-1MV 0V) (1MV, 10V) 
RCOMP	3	0	1MEG
*
* PWM OUTPUT STAGE
VCC	10	0	DC 10V
Q1	10	3 11	QNOM
RL1	11	0	20
*
* LINEAR OUTPUT STAGE
Q2	10	1 12	QNOM
RL2	12	0	20
*
.model	QNOM	NPN
*
* ANALYSIS
.TRAN 	5US  	2000US
* VIEW RESULTS
.PRINT	TRAN	V(1) V(3)
* TOPSPICE CALCULATIONS
*#CALC  PQ1=I(RL1)*(V(10)-V(11))
*#CALC  PQ2=I(RL2)*(V(10)-V(12))
.PROBE
.END
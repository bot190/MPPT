PWM_TRIAL_320
.LIB BRUTE_FORCE_VOLTAGE_SOURCE_320.LIB
.LIB BRUTE_FORCE_VOLTAGE_SOURCE_320_PERCENT.LIB
XV1 1 0 PWM
XV2 2 0 PERCENT
.PROBE
.TRAN 1580m 1580m 0u 1u UIC
.END